module vnoise
