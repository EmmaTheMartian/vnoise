module noise
